module sim_top();

timer_tb timer_test();
presc_tb presc_test();

endmodule
