module sim_top();

//timer_tb timer_test();
//presc_tb presc_test();
//spi_tb   spi_test();
//bcd_register_tb bcd_reg_test();
//ss_display_tb ss_display_test(); 
counter_tb counter_test();

endmodule
