module sim_top();

timer_tb timer_test();

endmodule
