// Nubmers in 7-segment encoding
`define SEG_0 7'b1111110
`define SEG_1 7'b0110000
`define SEG_2 7'b1101101
`define SEG_3 7'b1111001
`define SEG_4 7'b0110011
`define SEG_5 7'b1011011
`define SEG_6 7'b1011111
`define SEG_7 7'b1110000
`define SEG_8 7'b1111111
`define SEG_9 7'b1111011



