// Range of termperatures will vary from 0 to 100 degres of Celcius
module sim_top;
    //timer_tb timer_test();
    //presc_tb presc_test();
    register_tb register_test();
endmodule
