module sim_top();

endmodule
